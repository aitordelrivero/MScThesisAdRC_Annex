"SingleStageCascode"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Restart\cir\SingleStageCascode.asc
R3 N002 0 {Rs}
R4 N002 N003 {Ree}
C3 N002 N003 {Ce}
G1 0 N003 out 0 {1/gain}
I1 N002 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
XU1 N001 N003 0 0 CMOS18N W={W} L={L} ID={ID}
XU2 out 0 N001 N001 CMOS18N W={W} L={L} ID={ID}
.lib SLiCAP.lib
* W?
* loop reference?
.backanno
.end
