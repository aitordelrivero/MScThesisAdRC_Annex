mosEKVplots
* SLiCAP netlist file
.include SLiCAP.lib
X1 d g s 0 CMOS18N_V W={W} L={L} VD={V_D} VG={V_G} VS={V_S}
.param V_D=1.65 V_G=1.2 V_S=0 W=1u L=350n
.end
