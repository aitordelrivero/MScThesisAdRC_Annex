"CIRCUIT3IC"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\CIRCUIT3IC.asc
R3 N003 0 {Rs}
R4 N003 N001 {Ree}
C3 N003 N001 {Ce}
I1 N003 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
R1 N001 out {gain}
XU1 N002 out N001 0 CMOS18NDIC IC={ICas} L={Lin} ID={IDas}
XU2 N002 N002 0 0 CMOS18NIC IC={ICcm} L={Lcm} ID={IDasPMOS}
XU3 out N002 0 0 CMOS18NIC IC={ICcm} L={Lcm} ID={IDasPMOS}
.lib SLiCAP.lib
* loopgain reference: Gm_M1_XU1 (cascoded version, no Cdg)
* -
* -
* +
* +
* -
.backanno
.end
