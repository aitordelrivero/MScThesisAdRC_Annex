"LikelySelection"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\LikelySelection.asc
R3 N003 0 {Rs}
R4 N003 N001 {Ree}
C3 N003 N001 {Ce}
I1 N003 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
XU1 out N002 0 0 CMOS18N W={Wout} L={L} ID={IDout}
R1 N001 out {gain}
XU2 NC_01 N002 N001 0 CMOS18ND W={Was} L={L} ID={IDas}
.lib SLiCAP.lib
* loopgain reference: Gm_M1_XU1 (cascoded version, no Cdg)
* +
* +
* -
* -
* +
* +
* -
* -
* -
.backanno
.end
