"NoiseControllerAndFeedbackPMOS"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\NoiseControllerAndFeedbackPMOS.asc
XU1 N002 0 N003 PM18_noise ID={ID} IG={IG} W={W} L={L}
H1 out 0 N003 0 {gain}
R3 N001 0 {Rs}
R4 N001 N002 {Ree}
C3 N001 N002 {Ce}
In2 0 N002 I value=0 dc=0 dcvar=0 noise={4*k*T/gain}
R1 N002 0 {gain}
.lib SLiCAP.lib
.backanno
.end
