"DoubleStageVersion1"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\DoubleStageVersion1.asc
R3 N003 0 {Rs}
R4 N003 N001 {Ree}
C3 N003 N001 {Ce}
I1 N003 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
XU1 0 N002 out out CMOS18P W={Wout} L={Lout} ID={IDout}
R1 N001 out {gain}
XU2 0 N002 N001 0 CMOS18ND W={Was} L={Lin} ID={IDas}
.lib SLiCAP.lib
* loopgain reference: Gm_M1_XU2 (cascoded version, no Cdg)
* +
* +
* -
* -
* -
* -
* -
.backanno
.end
