"NoiseTIA"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\NoiseTIA.asc
In2 0 N002 I value=0 dc=0 dcvar=0 noise={4*k*T/gain}
R4 N001 0 {Rs}
R5 N001 N002 {Ree}
C3 N001 N002 {Ce}
In1 N002 N001 I value=0 dc=0 dcvar=0 noise={4*k*T/Ree}
In3 N001 0 I value=0 dc=0 dcvar=0 noise={4*k*T/Rs}
XU1 N002 0 N003 NM18_noise ID={ID} IG={IG} W={W} L={L}
H1 out 0 N003 0 {gain}
R1 N002 0 {gain}
.lib SLiCAP.lib
.backanno
.end
