"DoubleCSIdeal"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\DoubleCSIdeal.asc
R3 N003 0 {Rs}
R4 N003 N001 {Ree}
C3 N003 N001 {Ce}
I1 N003 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
XU1 N002 N001 0 0 CMOS18N W={W} L={L} ID={ID}
XU2 out P001 0 0 CMOS18N W={Wout} L={L} ID={IDout}
F1 P001 0 N002 0 1
R1 N001 out {gain}
.lib SLiCAP.lib
.backanno
.end
