"CIRCUIT6"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\AlternativeTopology\cir\CIRCUIT6.asc
R3 N004 0 {Rs}
R4 N004 N003 {Ree}
C3 N004 N003 {Ce}
I1 N004 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
R1 N003 out {gain}
XU1 N001 N002 N003 0 CMOS18ND W={Was} L={Lin} ID={IDas}
XU2 N001 N001 0 0 CMOS18P W={Wcm} L={Lcm} ID={IDasPMOS}
XU3 N002 N001 0 0 CMOS18P W={Wcm} L={Lcm} ID={IDasPMOS}
XU4 out N002 0 0 CMOS18P W={Wout} L={Lout} ID={IDoutPMOS}
XU5 out 0 0 0 CMOS18N W={Wb} L={Lb} ID={IDout}
XU6 NC_01 0 0 0 CMOS18N W={Wbcm} L={Lbcm} ID={2*IDas}
.lib SLiCAP.lib
* +
* -
* -
* -
.backanno
.end
