"FreqComp_Phantom_NoBias"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\New\cir\FreqComp_Phantom_NoBias.asc
R3 N004 0 {Rs}
R4 N004 N003 {Ree}
C3 N004 N003 {Ce}
I1 N004 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
R1 N003 N002 {gain}
XU1 0 N001 N003 0 CMOS18ND W={Was} L={Lin} ID={IDas}
XU4 N002 N001 0 0 CMOS18P W={Wout} L={Lout} ID={IDoutPMOS}
R2 N002 out {Rph1}
.lib SLiCAP.lib
* +
* -
* -
.backanno
.end
