"CIRCUIT2IC"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Passive\cir\CIRCUIT2IC.asc
R3 N002 0 {Rs}
R4 N002 N001 {Ree}
C3 N002 N001 {Ce}
I1 N002 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
R1 N001 out {gain}
XU1 0 out N001 0 CMOS18NDIC IC={ICas} L={Lin} ID={IDas}
.lib SLiCAP.lib
* loopgain reference: Gm_M1_XU1 (cascoded version, no Cdg)
* +
* -
* -
.backanno
.end
