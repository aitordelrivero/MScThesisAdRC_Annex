"CIRCUIT2"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\AlternativeTopology\cir\CIRCUIT2.asc
R3 N002 0 {Rs}
R4 N002 N001 {Ree}
C3 N002 N001 {Ce}
I1 N002 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
R1 N001 out {gain}
XU1 out 0 N001 0 CMOS18ND W={Was} L={Lin} ID={IDas}
.lib SLiCAP.lib
* +
* -
* -
.backanno
.end
