"DoubleCS"
* C:\Users\aitor\OneDrive\Msc Thesis\Chap2 Voltage clamp\Restart\cir\DoubleCS.asc
R3 N003 0 {Rs}
R4 N003 N004 {Ree}
C3 N003 N004 {Ce}
G1 0 N004 out 0 {1/gain}
I1 N003 0 I value=0 dc=0 dcvar=0 noise=0
C1 out 0 {Cload}
XU1 N001 N004 0 0 CMOS18N W={W} L={L} ID={ID}
XU2 out N002 0 0 CMOS18N W={Wout} L={L} ID={IDout}
XU3 N002 N001 0 0 CMOS18P W={Wcurmir} L={L} ID={ID}
XU4 N001 N001 0 0 CMOS18P W={Wcurmir} L={L} ID={ID}
.lib SLiCAP.lib
* PMOS CURRENT MIRROR to introduce a -1: \n- Use a low transconductance\n- Use a high cut-off frequency\n- Introduces a pole around ft/2
.backanno
.end
